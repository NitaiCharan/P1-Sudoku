�]q (]q(]q(]q(}q(X   digitoqX   5qX
   automaticoq�u}q(hX   4q	h�u}q
(hX   3qh�ue]q(}q(hX   8qh�u}q(hX   7qh�u}q(hX   6qh�ue]q(}q(hX   2qh�u}q(hX   1qh�u}q(hX   9qh�uee]q(]q(}q(hhh�u}q(hhh�u}q(hhh�ue]q(}q (hhh�u}q!(hhh�u}q"(hhh�ue]q#(}q$(hhh�u}q%(hhh�u}q&(hh	h�uee]q'(]q((}q)(hhh�u}q*(hhh�u}q+(hhh�ue]q,(}q-(hh	h�u}q.(hhh�u}q/(hhh�ue]q0(}q1(hhh�u}q2(hhh�u}q3(hhh�ueee]q4(]q5(]q6(}q7(hhh�u}q8(hhh�u}q9(hhh�ue]q:(}q;(hhh�u}q<(hhh�u}q=(hhh�ue]q>(}q?(hh	h�u}q@(hhh�u}qA(hhh�uee]qB(]qC(}qD(hhh�u}qE(hhh�u}qF(hhh�ue]qG(}qH(hh	h�u}qI(hhh�u}qJ(hhh�ue]qK(}qL(hhh�u}qM(hhh�u}qN(hhh�uee]qO(]qP(}qQ(hhh�u}qR(hhh�u}qS(hh	h�ue]qT(}qU(hhh�u}qV(hhh�u}qW(hhh�ue]qX(}qY(hhh�u}qZ(hhh�u}q[(hhh�ueee]q\(]q](]q^(}q_(hhh�u}q`(hhh�u}qa(hhh�ue]qb(}qc(hhh�u}qd(hhh�u}qe(hh	h�ue]qf(}qg(hhh�u}qh(hhh�u}qi(hhh�uee]qj(]qk(}ql(hhh�u}qm(hhh�u}qn(hhh�ue]qo(}qp(hhh�u}qq(hhh�u}qr(hhh�ue]qs(}qt(hhh�u}qu(hh	h�u}qv(hhh�uee]qw(]qx(}qy(hhh�u}qz(hh	h�u}q{(hhh�ue]q|(}q}(hhh�u}q~(hhh�u}q(hhh�ue]q�(}q�(hhh�u}q�(hhh�u}q�(hhh�ueeee.