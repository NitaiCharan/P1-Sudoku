�]q (]q(]q(]q(}q(X   digitoqX   5qX
   automaticoq�u}q(hX   4q	h�u}q
(hX   3qh�ue]q(}q(hX   1qh�u}q(hhh�u}q(hX   6qh�ue]q(}q(hhh�u}q(hhh�u}q(hX   9qh�uee]q(]q(}q(hhh�u}q(hhh�u}q(hhh�ue]q(}q(hX   2qh�u}q(hhh�u}q (hhh�ue]q!(}q"(hhh�u}q#(hhh�u}q$(hhh�uee]q%(]q&(}q'(hhh�u}q((hhh�u}q)(hhh�ue]q*(}q+(hh	h�u}q,(hhh�u}q-(hhh�ue]q.(}q/(hX   7q0h�u}q1(hhh�u}q2(hhh�ueee]q3(]q4(]q5(}q6(hhh�u}q7(hhh�u}q8(hhh�ue]q9(}q:(hhh�u}q;(hhh�u}q<(hhh�ue]q=(}q>(hhh�u}q?(hhh�u}q@(hhh�uee]qA(]qB(}qC(hhh�u}qD(hhh�u}qE(hhh�ue]qF(}qG(hh	h�u}qH(hhh�u}qI(hhh�ue]qJ(}qK(hhh�u}qL(hhh�u}qM(hhh�uee]qN(]qO(}qP(hhh�u}qQ(hhh�u}qR(hhh�ue]qS(}qT(hhh�u}qU(hhh�u}qV(hh0h�ue]qW(}qX(hhh�u}qY(hhh�u}qZ(hhh�ueee]q[(]q\(]q](}q^(hhh�u}q_(hX   8q`h�u}qa(hh0h�ue]qb(}qc(hhh�u}qd(hhh�u}qe(hh	h�ue]qf(}qg(hhh�u}qh(hhh�u}qi(hhh�uee]qj(]qk(}ql(hhh�u}qm(hhh�u}qn(hhh�ue]qo(}qp(hhh�u}qq(hhh�u}qr(hh`h�ue]qs(}qt(hhh�u}qu(hh	h�u}qv(hhh�uee]qw(]qx(}qy(hhh�u}qz(hh	h�u}q{(hhh�ue]q|(}q}(hhh�u}q~(hhh�u}q(hhh�ue]q�(}q�(hh`h�u}q�(hh0h�u}q�(hhh�ueeee.